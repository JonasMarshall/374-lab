//module ALU (input [31:0] A, B, input [3:0] op_sel, output [31:0] C);
//	begin 
//	end
// endmodule